module Top();
    frequency f1(JA, clk, an, seg);

endmodule