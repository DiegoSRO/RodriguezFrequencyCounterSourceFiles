module top()
        frequency f1(JA, clk, an, seg);
 //was not able to implement, JA is PMOD, clk is system clock, an is anode number that controls digit, seg is segment pattern
 //Cannot test this
endmodule